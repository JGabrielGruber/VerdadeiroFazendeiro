module models

import models { Producao, Terreno }

pub struct Plantio {
	producao Producao
	terreno Terreno
}
