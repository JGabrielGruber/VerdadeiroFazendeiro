module models

struct Proprietario {
	uid string
	mut:
		nome string
}
