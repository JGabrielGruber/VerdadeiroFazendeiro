module main

import src { run }

fn main() {
	println('Hello World!')
	run()
}
