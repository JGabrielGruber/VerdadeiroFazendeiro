module models

import models { Producao, Terreno }

struct Plantio {
	producao Producao
	terreno Terreno
}
