module models

pub struct Proprietario {
	uid string
	mut:
		nome string
}
