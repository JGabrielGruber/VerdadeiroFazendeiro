module models

pub struct Cultura {
	nome string
	tempo i64
	peso int // gramas
	mut:
		valor i64 // centavos
}
